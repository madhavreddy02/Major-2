
`timescale 1ns / 1ps

module mult_block #(IMAGE_SIZE = 16, KERNEL_SIZE = 3,EXP_SIZE = 5, MANT_SIZE = 10, DATA_WIDTH=8, ADDR_SIZE=4,MAX_ADDRESS=15, COLUMNS = 4, ROWS = 3)
(
input      [MANT_SIZE:0] I1, I2, I3, I4, I5, I6, I7, I8, I9,
input      [MANT_SIZE:0] K1, K2, K3, K4, K5, K6, K7, K8, K9,
output reg [(2 * MANT_SIZE):0] sign_mant_p1, sign_mant_p2, sign_mant_p3, sign_mant_p4, sign_mant_p5,
                               sign_mant_p6, sign_mant_p7, sign_mant_p8, sign_mant_p9         
);


multiplier #(.IMAGE_SIZE(IMAGE_SIZE), .KERNEL_SIZE(KERNEL_SIZE),.EXP_SIZE(EXP_SIZE) , .MANT_SIZE(MANT_SIZE) , .DATA_WIDTH(DATA_WIDTH), .ADDR_SIZE(ADDR_SIZE), .MAX_ADDRESS(MAX_ADDRESS), .COLUMNS(COLUMNS), .ROWS(ROWS)) M1 (.I(I1),.K(K1),.sign_mant_p(sign_mant_p1));
multiplier #(.IMAGE_SIZE(IMAGE_SIZE), .KERNEL_SIZE(KERNEL_SIZE),.EXP_SIZE(EXP_SIZE) , .MANT_SIZE(MANT_SIZE) , .DATA_WIDTH(DATA_WIDTH), .ADDR_SIZE(ADDR_SIZE), .MAX_ADDRESS(MAX_ADDRESS), .COLUMNS(COLUMNS), .ROWS(ROWS)) M2 (.I(I2),.K(K2),.sign_mant_p(sign_mant_p2));
multiplier #(.IMAGE_SIZE(IMAGE_SIZE), .KERNEL_SIZE(KERNEL_SIZE),.EXP_SIZE(EXP_SIZE) , .MANT_SIZE(MANT_SIZE) , .DATA_WIDTH(DATA_WIDTH), .ADDR_SIZE(ADDR_SIZE), .MAX_ADDRESS(MAX_ADDRESS), .COLUMNS(COLUMNS), .ROWS(ROWS)) M3 (.I(I3),.K(K3),.sign_mant_p(sign_mant_p3));
multiplier #(.IMAGE_SIZE(IMAGE_SIZE), .KERNEL_SIZE(KERNEL_SIZE),.EXP_SIZE(EXP_SIZE) , .MANT_SIZE(MANT_SIZE) , .DATA_WIDTH(DATA_WIDTH), .ADDR_SIZE(ADDR_SIZE), .MAX_ADDRESS(MAX_ADDRESS), .COLUMNS(COLUMNS), .ROWS(ROWS)) M4 (.I(I4),.K(K4),.sign_mant_p(sign_mant_p4));
multiplier #(.IMAGE_SIZE(IMAGE_SIZE), .KERNEL_SIZE(KERNEL_SIZE),.EXP_SIZE(EXP_SIZE) , .MANT_SIZE(MANT_SIZE) , .DATA_WIDTH(DATA_WIDTH), .ADDR_SIZE(ADDR_SIZE), .MAX_ADDRESS(MAX_ADDRESS), .COLUMNS(COLUMNS), .ROWS(ROWS)) M5 (.I(I5),.K(K5),.sign_mant_p(sign_mant_p5));
multiplier #(.IMAGE_SIZE(IMAGE_SIZE), .KERNEL_SIZE(KERNEL_SIZE),.EXP_SIZE(EXP_SIZE) , .MANT_SIZE(MANT_SIZE) , .DATA_WIDTH(DATA_WIDTH), .ADDR_SIZE(ADDR_SIZE), .MAX_ADDRESS(MAX_ADDRESS), .COLUMNS(COLUMNS), .ROWS(ROWS)) M6 (.I(I6),.K(K6),.sign_mant_p(sign_mant_p6));
multiplier #(.IMAGE_SIZE(IMAGE_SIZE), .KERNEL_SIZE(KERNEL_SIZE),.EXP_SIZE(EXP_SIZE) , .MANT_SIZE(MANT_SIZE) , .DATA_WIDTH(DATA_WIDTH), .ADDR_SIZE(ADDR_SIZE), .MAX_ADDRESS(MAX_ADDRESS), .COLUMNS(COLUMNS), .ROWS(ROWS)) M7 (.I(I7),.K(K7),.sign_mant_p(sign_mant_p7));
multiplier #(.IMAGE_SIZE(IMAGE_SIZE), .KERNEL_SIZE(KERNEL_SIZE),.EXP_SIZE(EXP_SIZE) , .MANT_SIZE(MANT_SIZE) , .DATA_WIDTH(DATA_WIDTH), .ADDR_SIZE(ADDR_SIZE), .MAX_ADDRESS(MAX_ADDRESS), .COLUMNS(COLUMNS), .ROWS(ROWS)) M8 (.I(I8),.K(K8),.sign_mant_p(sign_mant_p8));
multiplier #(.IMAGE_SIZE(IMAGE_SIZE), .KERNEL_SIZE(KERNEL_SIZE),.EXP_SIZE(EXP_SIZE) , .MANT_SIZE(MANT_SIZE) , .DATA_WIDTH(DATA_WIDTH), .ADDR_SIZE(ADDR_SIZE), .MAX_ADDRESS(MAX_ADDRESS), .COLUMNS(COLUMNS), .ROWS(ROWS)) M9 (.I(I9),.K(K9),.sign_mant_p(sign_mant_p9));

endmodule








